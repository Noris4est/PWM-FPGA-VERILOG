`timescale 1ns/1ps
module PWM_FPGA_TB1
#(
	parameter CLOCK_FREQUENCY			=400000,
	parameter PWM_FREQUENCY				=100000,
	parameter MAX_VALUE					=4,
	parameter DEEP_FILL_FACTOR			=$clog2(MAX_VALUE)+1
);
localparam PERIOD_IN_CLOCK_NS=1000000000/CLOCK_FREQUENCY;

reg	IN_CLOCK,IN_RESET,IN_ENABLE;
reg	[DEEP_FILL_FACTOR-1:0] 	IN_FILL_FACTOR;
wire OUT_PWM_SIGNAL;


PWM_FPGA
#(
	.CLOCK_FREQUENCY(CLOCK_FREQUENCY),
	.PWM_FREQUENCY(PWM_FREQUENCY),
	.MAX_VALUE(MAX_VALUE)
)
PWM_MODULE
(
	IN_CLOCK,
	IN_RESET,
	IN_ENABLE,
	IN_FILL_FACTOR,
	OUT_PWM_SIGNAL
);

initial begin
	IN_CLOCK=0;
	IN_RESET=0;
	IN_ENABLE=0;
end
always 
	begin
		#(PERIOD_IN_CLOCK_NS/2)
		IN_CLOCK=!IN_CLOCK;
	end
	
	
initial begin
	#(PERIOD_IN_CLOCK_NS*10)
	IN_FILL_FACTOR=2;	
	#(PERIOD_IN_CLOCK_NS*3)
	IN_RESET=1;
	#(PERIOD_IN_CLOCK_NS*8)
	IN_RESET=0;
	#(PERIOD_IN_CLOCK_NS*12)
	IN_ENABLE=1;
	#(PERIOD_IN_CLOCK_NS*30)
	IN_FILL_FACTOR=3;	
	#(PERIOD_IN_CLOCK_NS*5)
	IN_RESET=1;
	#(PERIOD_IN_CLOCK_NS*40)
	IN_RESET=0;
	#(PERIOD_IN_CLOCK_NS*3)
	IN_FILL_FACTOR=1;	
	#(PERIOD_IN_CLOCK_NS*2)
	IN_RESET=1;
	#(PERIOD_IN_CLOCK_NS*3)
	IN_RESET=0;
	#(PERIOD_IN_CLOCK_NS*30)
	IN_FILL_FACTOR=0;
	#(PERIOD_IN_CLOCK_NS*3)
	IN_RESET=1;
	#(PERIOD_IN_CLOCK_NS*3)
	IN_RESET=0;
	#(PERIOD_IN_CLOCK_NS*30)
	IN_FILL_FACTOR=4;
	#(PERIOD_IN_CLOCK_NS*3)
	IN_RESET=1;
	#(PERIOD_IN_CLOCK_NS*3)
	IN_RESET=0;
end

endmodule
